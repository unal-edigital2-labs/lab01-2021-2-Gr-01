`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:26:57 08/19/2019 
// Design Name: 
// Module Name:    sum1bcc 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////

module sum1bcc (A, B, Ci, Cout, S);

  input  wire A;
  input  wire B;
  input  wire Ci;
  output wire Cout;
  output wire S;

  wire [1:0] st;
  assign S = st[0];
  assign Cout = st[1];

  assign st = A + B + Ci;
 
  
endmodule

